<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML+RDFa 1.0//EN" "http://www.w3.org/MarkUp/DTD/xhtml-rdfa-1.dtd">
<html xmlns="http://www.w3.org/1999/xhtml" xmlns:cc="http://creativecommons.org/ns#" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:dct="http://purl.org/dc/terms/" xmlns:frbr="http://purl.org/vocab/frbr/core#" xml:lang="sv">
<head about="http://creativecommons.org/licenses/by-sa/3.0/">
<meta name="viewport" content="width=device-width, initial-scale=1.0" />
<meta http-equiv="Content-Type" content="application/xhtml+xml; charset=utf-8" />
<title>Creative Commons &mdash; Erkännande-DelaLika 3.0 Unported
  &mdash; CC BY-SA 3.0 </title>
<meta http-equiv="content-type" content="text/html;charset=utf-8" />
<link rel="stylesheet" href="//maxcdn.bootstrapcdn.com/bootstrap/3.3.7/css/bootstrap.min.css" integrity="sha384-BVYiiSIFeK1dGmJRAkycuHAHRg32OmUcww7on3RYdg4Va+PmSTsz/K68vbdEjh4u" crossorigin="anonymous">
<link rel='stylesheet' id='cc-google-fonts-css' href='//fonts.googleapis.com/css?family=Source+Sans+Pro%3A400%2C600%2C700%7CRoboto+Condensed' type='text/css' media='all' />
<link rel='stylesheet' id='cc-fontello-css' href="/wp-content/themes/cc/fonts/fontello/css/cc-fontello.css" type='text/css' media='all' />
<link rel="stylesheet" id="twentysixteen-jetpack-css" href="/wp-content/plugins/jetpack/modules/theme-tools/compat/twentysixteen.css" type="text/css" media="all">
<link rel='stylesheet' id='parent-style-css' href="/wp-content/themes/twentysixteen/style.css" type='text/css' media='all' />
<link rel='stylesheet' id='cc-style-css' href="/wp-content/themes/cc/css/app.css" type='text/css' media='all' />
<link rel="stylesheet" type="text/css" href="/includes/deed4.css" media="screen" />
<link rel="stylesheet" type="text/css" media="print" href="/includes/deed4-print.css" />
<link rel="stylesheet" type="text/css" href="/includes/jurisdictions.css" media="screen" />
<!--[if lt IE 7]>
    <link rel="stylesheet" type="text/css"
          href="/includes/deed3-ie.css"
          media="screen" />
  <![endif]-->
<link rel="alternate" type="application/rdf+xml" href="rdf" />
<script type="text/javascript">
function setCookie(name, value, expires, path, domain, secure) {
    document.cookie= name + "=" + escape(value) +
        ((expires) ? "; expires=" + expires.toGMTString() : "") +
        ((path) ? "; path=" + path : "") +
        ((domain) ? "; domain=" + domain : "") +
        ((secure) ? "; secure" : "");
}
var expiry = new Date();
expiry.setTime(expiry.getTime()+(5*365*24*60*60*1000));
setCookie('lang','%s', expiry, '/');
</script>
<script src="https://cdnjs.cloudflare.com/ajax/libs/tether/1.4.0/js/tether.min.js"></script>
<script src="https://cdnjs.cloudflare.com/ajax/libs/jquery/1.12.4/jquery.min.js" integrity="sha384-nvAa0+6Qg9clwYCGGPpDQLVpLNn0fRaROjHqs13t4Ggj3Ez50XnGQqc/r8MhnRDZ" crossorigin="anonymous"></script>
<script src="https://maxcdn.bootstrapcdn.com/bootstrap/3.3.7/js/bootstrap.min.js" integrity="sha384-Tc5IQib027qvyjSMfHjOMaLkfuWVxZxUPnCJA7l2mCWNIpG9mGCD8wGNIcPD7Txa" crossorigin="anonymous"></script>
</head>
<body typeof="cc:License" about="http://creativecommons.org/licenses/by/4.0/" class="license ltr">


<div id="page" class="site">
<div class="site-inner">
<a class="skip-link screen-reader-text" href="#content">Hoppa över till innehåll</a>
<div class="site-header-wrapper">
<header id="masthead" class="site-header sticky-nav-main" role="banner">
<div class="site-header-main">
<div class="site-branding">
<a class="cc-site-logo-link" href="https://creativecommons.org/" rel="home">
<img class="cc-site-logo" width="303" height="72" src="https://creativecommons.org/wp-content/themes/cc/images/cc.logo.white.svg">
</a>
</div>
<button id="menu-toggle" class="menu-toggle"><i class="cc-icon-menu"></i> <span>Meny</span></button>
<div id="site-header-menu" class="site-header-menu">
<nav id="mobile-navigation" class="mobile-navigation" role="navigation" aria-label="Mobile Menu">
<div class="menu-mobile-menu-container"><ul id="menu-mobile-menu" class="mobile-menu">
<li id="menu-item-48798" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48798"><a href="https://creativecommons.org/share-your-work/">Dela ditt arbete</a></li>
<li id="menu-item-48799" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48799"><a href="https://creativecommons.org/use-remix/">Använd &#038; remix</a></li>
<li id="menu-item-48800" class="menu-item menu-item-type-post_type menu-item-object-page page_item page-item-7466 menu-item-48800"><a href="https://creativecommons.org/about/">What We do</a></li>
<li id="menu-item-48801" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48801"><a href="https://creativecommons.org/blog/">Blogg</a></li>
<li id="menu-item-48802" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48802"><a href="https://network.creativecommons.org/?ref=global-affiliate-network">Global Network</a></li>
<li id="menu-item-48803" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48803"><a href="https://creativecommons.org/use-remix/search-the-commons/">Sök i Commons</a></li>
</ul></div>
</nav>
<nav id="site-navigation" class="main-navigation" role="navigation" aria-label="Primary Menu">
<div class="menu-primary-menu-container"><ul id="menu-primary-menu" class="primary-menu">
<li id="menu-item-48791" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48791"><a href="https://creativecommons.org/share-your-work/">Dela ditt arbete</a></li>
<li id="menu-item-48792" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48792"><a href="https://creativecommons.org/use-remix/">Använd &#038; remix</a></li>
<li id="menu-item-48570" class="menu-item menu-item-type-post_type menu-item-object-page page_item page-item-7466 menu-item-48570"><a href="https://creativecommons.org/about/">What We do</a></li>
<li id="menu-item-48793" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48793"><a href="https://creativecommons.org/blog/">Blogg</a></li>
</ul></div>
</nav>
<nav id="secondary-navigation" class="secondary-navigation" role="navigation" aria-label="Secondary Menu">
<div class="menu-secondary-menu-container"><ul id="menu-secondary-menu" class="secondary-menu">
<li id="menu-item-55890" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-55890"><a href="https://search.creativecommons.org/">Search for CC images</a></li>
<li id="menu-item-48804" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48804"><a href="https://network.creativecommons.org/?ref=global-affiliate-network">Global Network</a></li>
<li id="menu-item-56460" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-56460"><a href="https://us.e-activist.com/page/6747/subscribe/1?ea.tracking.id=mailing-list-page">Newsletters</a></li>
<li id="menu-item-52800" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-52800"><a href="https://store.creativecommons.org/">Store</a></li>
<li id="menu-item-48806" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48806"><a href="https://creativecommons.org/about/contact/">Kontakt</a></li>
</ul></div>
</nav>
<nav id="social-navigation" class="social-navigation" role="navigation" aria-label="Social Links Menu">
<div class="menu-social-links-container"><ul id="menu-social-links" class="social-links-menu">
<li id="menu-item-48807" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48807"><a href="https://www.facebook.com/creativecommons"><span class="screen-reader-text">Facebook</span></a></li>
<li id="menu-item-48808" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48808"><a href="https://twitter.com/creativecommons"><span class="screen-reader-text">Twitter</span></a></li>
<li id="menu-item-48809" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-48809"><a href="mailto:info@creativecommons.org"><span class="screen-reader-text">E-post</span></a></li>
</ul></div>
</nav>
</div>
</div>
</header>
</div>
<div id="content" class="site-content">
<aside id="header-below" class="widget-area">
<section id="text-15" class="widget-1 widget-first widget-last widget-odd widget widget_text">
<div class="textwidget">
<div id="donation-bar-wrapper" class="donation-bar-wrapper">
<div id="donation-bar-inner" class="donation-bar-inner">
<p class="donate-text">Hjälp oss bygga ett livfullt, globalt sammarbetande commons</p>
<div class="donate-action"><a href="https://us.netdonor.net/page/6650/donate/1?ea.tracking.id=deed-top" class="button donate arrow">Donera<span class="hide-on-mobile"> Nu</span></a></div>
</div>
</div>
</div>
</section>
</aside>
<div id="language-selector-block" class="container">
<div class="language-selector-inner">
<span dir="ltr" style="text-align: left">
Denna sida finns tillgänglig på följande språk:
</span>
<img class="language-icon" src="/images/language_icon_x2.png" alt="Languages" />
<select>
<option value="id">
Bahasa Indonesia
</option>
<option value="ms">
Bahasa Malaysia
</option>
<option value="es_ES">
Castellano (España)
</option>
<option value="ca">
Català
</option>
<option value="da">
Dansk
</option>
<option value="de">
Deutsch
</option>
<option value="en">
English
</option>
<option value="es">
Español
</option>
<option value="eo">
Esperanto
</option>
<option value="eu">
Euskara
</option>
<option value="fr">
français
</option>
<option value="gl">
Galego
</option>
<option value="hr">
hrvatski
</option>
<option value="it">
Italiano
</option>
<option value="lv">
Latviski
</option>
<option value="lt">
Lietuvių
</option>
<option value="hu">
Magyar
</option>
<option value="nl">
Nederlands
</option>
<option value="no">
norsk
</option>
<option value="pl">
polski
</option>
<option value="pt">
Português
</option>
<option value="pt_BR">
Português (BR)
</option>
<option value="ro">
română
</option>
<option value="sl">
Slovenščina
</option>
<option value="sr_LATN">
srpski (latinica)
</option>
 <option value="fi">
suomeksi
</option>
<option value="sv" selected="selected">
svenska
</option>
<option value="tr">
Türkçe
</option>
<option value="is">
Íslenska
</option>
<option value="cs">
čeština
</option>
<option value="el">
Ελληνικά
</option>
<option value="be">
Беларуская
</option>
<option value="ru">
русский
</option>
<option value="uk">
українська
</option>
<option value="ar">
العربية
</option>
<option value="fa">
پارسی
</option>
<option value="bn">
বাংলা
</option>
<option value="zh">
中文
</option>
<option value="ja">
日本語
</option>
<option value="zh_TW">
華語 (台灣)
</option>
<option value="ko">
한국어
</option>
</select>
</div>
</div>
<div id="primary" class="content-area">
<main id="main" class="site-main container" role="main">
<div id="deed" class="row" dir="ltr" style="text-align: left">
<div id="deed-head" class="row">
<div class="print-only icon cc-logo-print">
<img alt="cc logo" src="/images/deed/cc-logo.jpg">
</div>
<div id="cc-link">
<a rel="dc:creator dct:creator" href="/">
<span property="dc:title dct:title">Creative Commons</span>
</a>
</div>
<h1><span>Creative Commons Licens Deed</span></h1>
<div id="deed-license">
<h2>
<span class="cc-license-icons">
<span id="cc-logo" class="icon"><img alt="cc logo" src="/images/deed/cc_icon_white_x2.png"></span>
<span id="cc-attribution" class="icon"><img src="/images/deed/attribution_icon_white_x2.png"></span>
<span id="cc-icon-sa" class="icon"><img src="/images/deed/sa_white_x2.png"></span>
</span>
<span class="cc-license-title" property="dc:title dct:title">Erkännande-DelaLika 3.0 Unported</span>
<span class="cc-license-identifier" property="dc:identifier dct:identifier">
(CC BY-SA 3.0)
</span>
</h2>
</div>
</div>
<div id="deed-main" dir="ltr" style="text-align: left" class="row">
<div id="legalcode-block">
<div id="deed-disclaimer">
<span class="summary">
Detta är en lättläst sammanfattning av (och inte en ersättning för) <a href="legalcode.sv" class="fulltext">licensen</a>.
</span>
<span class="disclaimer">
<a href="#" id="disclaimer_popup" class="helpLink">Friskrivning</a>.
</span>
</div>
</div>
<div id="deed-main-content" class="row ">
<div id="deed-rights" dir="ltr" style="text-align: left" class="row">
<div class="col-sm-offset-2 col-sm-8">
<h3 style="text-align: center" resource="http://creativecommons.org/ns#Reproduction" rel="cc:permits">Du har tillstånd att:</h3>
<ul class="license-properties">
<li class="license share" rel="cc:permits" resource="http://creativecommons.org/ns#Distribution">
<strong>Dela</strong> &mdash; kopiera och vidaredistribuera materialet oavsett medium eller format
</li>
<li class="license remix" rel="cc:permits" resource="http://creativecommons.org/ns#DerivativeWorks">
<strong>Bearbeta</strong> &mdash; remixa, transformera, och bygg vidare på materialet
</li>
<li class="license commercial">
för alla ändamål, även kommersiellt.
</li>
<li id="more-container" class="license-hidden">
<span id="devnations-container" />
</li>
</ul>
</div>
<div id="libre" class="col-sm-2">
<a href="https://freedomdefined.org/" class="screen-only">
<img src="/images/deed/FreeCulturalWorks_seal_x2.jpg" style="border: 0" alt="Med denna licens blir ditt verk " Fri kultur"." />
</a>
<a href="https://freedomdefined.org/" class="print-only">
<img src="/images/deed/seal.png" style="border: 0" alt="" />
</a>
</div>
</div>
<div class="row">
<ul id="license-freedoms-no-icons" style="text-align: center" class="col-sm-offset-2 col-sm-8">
<li class="license">Licensgivaren kan inte återkalla dessa friheter så länge du följer licensvillkoren.</li>
</ul>
</div>
<div class="row"><div class="col-md-offset-1 col-md-10"><hr /></div></div>
<div id="deed-conditions" class="row">
<h3 style="text-align: center">På följande villkor:</h3>
<ul dir="ltr" style="text-align: left" class="license-properties col-md-offset-2 col-md-8">
<li class="license by">
<p>
<strong>Erkännande</strong> &mdash; <span rel="cc:requires" resource="http://creativecommons.org/ns#Attribution">Du måste ge <a href="#" id="appropriate_credit_popup" class="helpLink">ett korrekt erkännande</a></span>, ange en hyperlänk till licensen, och <span rel="cc:requires" resource="http://creativecommons.org/ns#Notice"><a href="#" id="indicate_changes_popup" class="helpLink">ange om bearbetningar är gjorda </a></span>. Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att licensgivaren stödjer dig eller ditt användande.
<span id="by-more-container"></span>
</p>
<p id="work-attribution-container" style="display:none;">
<strong>
Erkänn detta arbete:
</strong>
<br />
<input id="work-attribution" value="" type="text" readonly="readonly" onclick="this.select()" onfocus="document.getElementById('work-attribution').select();" />
<input id="license-code" type="hidden" value="CC BY-SA 3.0" />
<input id="license-url" type="hidden" value="http://creativecommons.org/licenses/by-sa/3.0/" />
<a href="" id="attribution_help" class="helpLink">
<img src="/images/information.png" alt="Information" />
</a>
</p>
</li>
<li class="license sa" rel="cc:requires" resource="http://creativecommons.org/ns#ShareAlike">
<p>
<strong>DelaLika</strong> &mdash; Om du remixar, transformerar eller bygger vidare på materialet måste du distribuera dina bidrag under <a href="#" id="same_license_popup" class="helpLink">samma licens</a> som originalet.
<span id="sa-more-container"></span>
</p>
</li>
</ul>
</div>
<div class="row">
<ul id="deed-conditions-no-icons" class="col-md-offset-2 col-md-8">
<li class="license">
<strong>Inga ytterligare begränsningar</strong> &mdash; Du får inte tillämpa lagliga begränsningar eller <a href="#" id="technological_measures_popup" class="helpLink">teknologiska metoder</a> som juridiskt begränsar andra från att gör något som licensen tillåter.
</li>
</ul>
</div>
<div class="row"><div class="col-md-offset-1 col-md-10"><hr /></div></div>
<div id="deed-understanding" class="row">
<h3 style="text-align: center">
Anmärkningar:
</h3>
<ul class="understanding license-properties col-md-offset-2 col-md-8">
<li class="license">
Du behöver inte följa licensvillkoren för de delar av materialet som finns i public domain eller där ditt användande är tillåtet av en tillämplig <a href="#" id="exception_or_limitation_popup" class="helpLink">undantag eller begränsning</a>.
</li>
<li class="license">
Inga garantier ges. Licensen ger eller ger dig inte alla de nödvändiga villkoren för ditt tänkta användande av verket. Till exempel, andra rättigheter som <a href="#" id="publicity_privacy_or_moral_rights_popup" class="helpLink">publicitet, integritetslagstiftning, eller ideella rättigheter </a> kan begränsa hur du kan använda verket.
</li>
</ul>
</div>
<span id="referrer-metadata-container" />
</div>
</div>
<div class="row" id="footer">
<p class="learn-more-cc">
<a href="https://wiki.creativecommons.org/FAQ">Lär dig mer</a> om CC-licensiering, eller <a id="get_this" href="/choose/results-one?license_code=by-sa&amp;amp;jurisdiction=&amp;amp;version=3.0&amp;amp;lang=sv">använd licensen</a> för ditt eget material.
</p>
<noscript>
                  <div id="deed-donate-footer">
                    <div class="footer-trigger">
                      <img src="/images/deed/cc_heart_x2.png" class="footer-logo" alt="" width="133" height="117" />
                      <div class="footer-trigger-content">
                        <p>Detta innehåll är fritt tillgängligt under enkla juridiska termer eftersom Creative Commons är en ideell förening som är beroende av donationer. Om du tycker om  detta innehåll, och tycker om att det är gratis för alla, då tycker vi att du ska fundera på att bidra med en donation till stöd för vårt arbete.</p>
                        <a href="https://us.netdonor.net/page/6650/donate/1?ea.tracking.id=license-footer"><button>Make a Donation</button></a>
                      </div>
                    </div>
                  </div>
                </noscript>
<div id="languages">
<span dir="ltr" style="text-align: left">
Denna sida finns tillgänglig på följande språk:
</span>
<br />
<a title="Bahasa Indonesia" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.id" hreflang="id" xml:lang="id">Bahasa Indonesia</a>
<a title="Bahasa Malaysia" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ms" hreflang="ms" xml:lang="ms">Bahasa Malaysia</a>
<a title="Castellano (España)" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.es_ES" hreflang="es_ES" xml:lang="es_ES">Castellano (España)</a>
<a title="Català" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ca" hreflang="ca" xml:lang="ca">Català</a>
<a title="Dansk" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.da" hreflang="da" xml:lang="da">Dansk</a>
<a title="Deutsch" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.de" hreflang="de" xml:lang="de">Deutsch</a>
<a title="English" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.en" hreflang="en" xml:lang="en">English</a>
<a title="Español" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.es" hreflang="es" xml:lang="es">Español</a>
<a title="Esperanto" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.eo" hreflang="eo" xml:lang="eo">Esperanto</a>
<a title="Euskara" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.eu" hreflang="eu" xml:lang="eu">Euskara</a>
<a title="français" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.fr" hreflang="fr" xml:lang="fr">français</a>
<a title="Galego" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.gl" hreflang="gl" xml:lang="gl">Galego</a>
<a title="hrvatski" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.hr" hreflang="hr" xml:lang="hr">hrvatski</a>
<a title="Italiano" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.it" hreflang="it" xml:lang="it">Italiano</a>
<a title="Latviski" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.lv" hreflang="lv" xml:lang="lv">Latviski</a>
<a title="Lietuvių" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.lt" hreflang="lt" xml:lang="lt">Lietuvių</a>
<a title="Magyar" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.hu" hreflang="hu" xml:lang="hu">Magyar</a>
<a title="Nederlands" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.nl" hreflang="nl" xml:lang="nl">Nederlands</a>
<a title="norsk" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.no" hreflang="no" xml:lang="no">norsk</a>
<a title="polski" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.pl" hreflang="pl" xml:lang="pl">polski</a>
<a title="Português" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.pt" hreflang="pt" xml:lang="pt">Português</a>
<a title="Português (BR)" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.pt_BR" hreflang="pt_BR" xml:lang="pt_BR">Português (BR)</a>
<a title="română" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ro" hreflang="ro" xml:lang="ro">română</a>
<a title="Slovenščina" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.sl" hreflang="sl" xml:lang="sl">Slovenščina</a>
<a title="srpski (latinica)" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.sr_LATN" hreflang="sr_LATN" xml:lang="sr_LATN">srpski (latinica)</a>
<a title="suomeksi" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.fi" hreflang="fi" xml:lang="fi">suomeksi</a>
<a title="svenska" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.sv" hreflang="sv" xml:lang="sv">svenska</a>
<a title="Türkçe" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.tr" hreflang="tr" xml:lang="tr">Türkçe</a>
<a title="Íslenska" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.is" hreflang="is" xml:lang="is">Íslenska</a>
<a title="čeština" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.cs" hreflang="cs" xml:lang="cs">čeština</a>
<a title="Ελληνικά" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.el" hreflang="el" xml:lang="el">Ελληνικά</a>
<a title="Беларуская" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.be" hreflang="be" xml:lang="be">Беларуская</a>
<a title="русский" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ru" hreflang="ru" xml:lang="ru">русский</a>
<a title="українська" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.uk" hreflang="uk" xml:lang="uk">українська</a>
<a title="العربية" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ar" hreflang="ar" xml:lang="ar">العربية</a>
<a title="پارسی" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.fa" hreflang="fa" xml:lang="fa">پارسی</a>
<a title="বাংলা" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.bn" hreflang="bn" xml:lang="bn">বাংলা</a>
<a title="中文" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.zh" hreflang="zh" xml:lang="zh">中文</a>
<a title="日本語" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ja" hreflang="ja" xml:lang="ja">日本語</a>
<a title="華語 (台灣)" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.zh_TW" hreflang="zh_TW" xml:lang="zh_TW">華語 (台灣)</a>
<a title="한국어" rel="alternate nofollow frbr:translation" rev="frbr:translationOf" href="./deed.ko" hreflang="ko" xml:lang="ko">한국어</a>
</div>
</div>
<div id="deed-donate-slide" style="display: none;">
<div class="slide-trigger">
<div class="slide-close"></div>
<img src="/images/deed/logo-cc-heart-white.png" class="slide-logo" alt="" width="100" height="88" />
<p class="desktop-only">Detta innehåll är fritt tillgängligt under enkla juridiska termer eftersom Creative Commons är en ideell förening som är beroende av donationer. Om du tycker om detta innehåll, och tycker om att det är gratis för alla, då tycker vi att du ska fundera på att bidra med en donation till stöd för vårt arbete.</p>
<p class="mobile-only">När du delar med dig så vinner alla.</p>
<div class="donate-box">
<div class="widget-inner">
<div class="gform_wrapper" id="gform_wrapper_10">
<form method="get" id="gform_10" action="https://us.netdonor.net/page/6650/donate/1" class="deed-donate-form">
<div id="field_10_1" class="gfield field_sublabel_below field_description_below">
<label class="gfield_label">Bidrag idag till Creative Commons</label>
<div class="ginput_container ginput_container_radio">
<ul class="gfield_radio" id="input_10_1">
<li class="gchoice_10_1_0">
<input name="transaction.donationAmt" type="radio" value="5" id="choice_10_1_0" tabindex="1">
<label for="choice_10_1_0" id="label_10_1_0">$5</label>
</li>
<li class="gchoice_10_1_1">
<input name="transaction.donationAmt" type="radio" value="15" checked="checked" id="choice_10_1_1" tabindex="2">
<label for="choice_10_1_1" id="label_10_1_1">$15</label>
</li>
<li class="gchoice_10_1_2">
<input name="transaction.donationAmt" type="radio" value="25" id="choice_10_1_2" tabindex="3">
<label for="choice_10_1_2" id="label_10_1_2">$25</label>
</li>
<li class="gchoice_10_1_3">
<input name="transaction.donationAmt" type="radio" value="50" id="choice_10_1_3" tabindex="4">
<label for="choice_10_1_3" id="label_10_1_3">$50</label>
</li>
<li class="gchoice_10_1_4">
<input name="transaction.donationAmt" type="radio" value="gf_other_choice" id="choice_10_1_4" tabindex="5" onfocus="$(this).next('input').focus();">
<input name="transaction.donationAmt.other" type="text" id="input_10_1_other" tabindex="5" style="max-width: 80%" placeholder="Summa" aria-label="Summa">
</li>
</ul>
<input type="hidden" name="type" value="One Time">
<input type="hidden" name="ea.tracking.id" value="deed-overlay">
<input type="submit" id="gform_submit_button_10" class="gform_button button" value="Donera nu!" tabindex="6">
</div>
</div>
</form>
</div>
</div>
</div>
</div>
</div>
</div>
</main>
</div>
</div>
<div class="site-footer-wrapper">
<footer id="colophon" class="site-footer sticky-nav-main" role="contentinfo">
<div class="cc-footer">
<div class="column cc-footer-main">
<div class="cc-footer-logo">
<a href="https://creativecommons.org/" class="custom-logo-link" rel="home" itemprop="url"><img width="980" height="240" src="https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_.png" class="custom-logo" alt="cc.logo.white" itemprop="logo" srcset="https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_.png 980w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-300x73.png 300w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-768x188.png 768w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-140x34.png 140w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-50x12.png 50w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-270x66.png 270w, https://creativecommons.org/wp-content/uploads/2016/06/cc.logo_.white_-245x60.png 245w" sizes="(max-width: 709px) 85vw, (max-width: 909px) 67vw, (max-width: 1362px) 62vw, 840px" /></a>
</div>
<div class="cc-footer-links">
<div class="menu-footer-links-container">
<ul id="menu-footer-links" class="menu">
<li id="menu-item-48794" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48794"><a href="https://creativecommons.org/about/contact/">Kontakt</a></li>
<li id="menu-item-48795" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48795"><a href="https://creativecommons.org/privacy/">Integritet</a></li>
<li id="menu-item-48796" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48796"><a href="https://creativecommons.org/policies/">Policyer</a></li>
<li id="menu-item-48797" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-48797"><a href="https://creativecommons.org/terms/">Villkor</a></li>
</ul>
</div>
</div>
</div>
<div class="column cc-footer-contact">
<h6><a href="https://creativecommons.org/about/contact">Vi blir jätteglada om du hör av dig!</a></h6>
<address>
Creative Commons<br />
PO Box 1866, Mountain View, CA 94042
</address>
<ul>
<li><a href="mailto:info@creativecommons.org" class="mail">info@creativecommons.org</a></li>
<li><a href="https://creativecommons.org/faq">Vanliga frågor</a></li>
</ul>
</div>
<div class="column cc-footer-license">
<div class="license-icons">
<a rel="license" href="https://creativecommons.org/licenses/by/4.0/" title="Creative Commons Attribution 4.0 International license">
<i class="cc-icon-cc"></i>
<i class="cc-icon-cc-by"></i>
</a>
</div>
<aside>
<div xmlns:cc="https://creativecommons.org/ns#" about="https://creativecommons.org">
<p>Except where otherwise <a class="subfoot" href="https://creativecommons.org/policies#license">noted</a>, content on this site is licensed under a <a class="subfoot" href="https://creativecommons.org/licenses/by/4.0/" rel="license">Creative Commons Attribution 4.0 International license</a>. <a class="subfoot" href="https://creativecommons.org/website-icons" target="blank">Icons</a> by The Noun Project.</p>
</div>
</aside>
</div>
</div>
</footer>
</div>
</div>
</div>
<div id="help-panels" style="display: none">
<div id="help_disclaimer_popup" class="help_panel">
<div class="hd">Friskrivning</div>
<div class="bd">
<p>Denna sammanfattning uppmärksammar enbart vissa av de viktigaste inslagen och villkoren från den faktiska licensen. Den är inte en licens och har inget juridiskt värde. Du bör noggrant gå igenom alla villkor i den faktiska licensen innan du använder det licensierade materialet.</p>
<p>Creative Commons är ingen advokatbyrå och tillhandahåller inga juridiska tjänster eller juridisk rådgivning. Distribution eller visning av, samt länkning till denna handling eller licensen som sammanfattas skapar ingen advokat-klient- eller annat förhållande.</p>
</div>
</div>
<div id="help_attribution_help" class="help_panel">
<div class="hd">
Vad betyder "Erkänna detta verk"?
</div>
<div class="bd">
<p>Sidan du kom från innehöll inbäddad licensmetadata, inklusive hur skaparen vill bli omnämnd vid återanvändning. Du kan använda HTML-koden här för att referera till verket. Då kommer även metadata att inkluderas på din sida så att andra också kan hitta ursprungsverket.</p>
</div>
</div>
<div id="help_mediation_and_arbitration_popup" class="help_panel">
<div class="bd">
<p>De tillämpliga medlingsreglerna kommer att bestämmas utifrån de upphovsrättsliga begränsningar som publiceras med verket, eller om inga då ska beslut fattas vid krav om medling. Om inget annat finns angivet i Copyrights noteringarna som kopplas till verket, kommer UNCITRAL medlingsregler att används vid medlingsbeslut.</p>
<p><a href="https://wiki.creativecommons.org/Intergovernmental_Organizations#What_should_I_know_before_I_use_a_work_licensed_under_the_IGO_3.0_ported_licenses.3F">Mer information</a>.</p>
</div>
</div>
<div id="help_appropriate_credit_popup" class="help_panel">
<div class="bd">
<p>Om det anges, måste du ange namnet på upphovsmannen och skriva ut villkoren för upphovsmannen, licensen, friskrivningsklausul och länka till verket. CC licenser före version 4.0 kräver också att du anger titeln på verket om det anges, och kan ha andra små skillnader </p>
<p><a href="https://wiki.creativecommons.org/License_Versions#Detailed_attribution_comparison_chart">Mer information</a>.</p>
</div>
</div>
<div id="help_indicate_changes_popup" class="help_panel">
<div class="bd">
<p>I 4.0, måste du indikera om du har modifierat materialet samt behålla indikeringar på tidigare modifieringar. I 3.0 och tidigare licensversioner krävs indikering av ändringar endast om du skapar en bearbetning.</p>
<p><a href="https://wiki.creativecommons.org/Best_practices_for_attribution#This_is_a_good_attribution_for_material_you_modified_slightly">Märkningsguide</a>.</p>
<p><a href="https://wiki.creativecommons.org/License_Versions#Modifications_and_adaptations_must_be_marked_as_such ">Mer information</a>.</p>
</div>
</div>
<div id="help_same_license_popup" class="help_panel">
<div class="bd">
<p>Du kan även använd en licens som listas som likvärdig på <a href="https://creativecommons.org/compatiblelicenses">https://creativecommons.org/compatiblelicenses</a></p>
<p><a href="https://wiki.creativecommons.org/FAQ#If_I_derive_or_adapt_material_offered_under_a_Creative_Commons_license.2C_which_CC_license.28s.29_can_I_use.3F">Mer information</a>.</p>
</div>
</div>
<div id="help_commercial_purposes_popup" class="help_panel">
<div class="bd">
<p>En kommersiell användning är en som främst är avsedd för kommersiell nytta eller monetär ersättning. </p>
<p><a href="https://wiki.creativecommons.org/Frequently_Asked_Questions#Does_my_use_violate_the_NonCommercial_clause_of_the_licenses.3F">Mer information</a>.</p>
</div>
</div>
<div id="help_some_kinds_of_mods_popup" class="help_panel">
<div class="bd">
<p>Att enbart ändra formatet skapar aldrig en bearbetning.</p>
<p><a href="https://wiki.creativecommons.org/Frequently_Asked_Questions#When_is_my_use_considered_an_adaptation.3F">Mer information</a>.</p>
</div>
</div>
<div id="help_technological_measures_popup" class="help_panel">
<div class="bd">
<p>Licensen förbjuder applikationer av effektiva teknologiska medel definierad med hänvisning till Artikel 11 i WIPO Copyright Treaty, WIPOs Upphovsrättsfördrag.</p>
<p><a href="https://wiki.creativecommons.org/License_Versions#Application_of_effective_technological_measures_by_users_of_CC-licensed_works_prohibited">Mer information</a>.</p>
</div>
</div>
<div id="help_exception_or_limitation_popup" class="help_panel">
<div class="bd">
<p>Rätten att använda verket enligt de undantag och begränsningar som finns i lagstiftningen, t.ex citaträtten, begränsas inte av CC licenserna. </p>
<p><a href="https://wiki.creativecommons.org/Frequently_Asked_Questions#Do_Creative_Commons_licenses_affect_exceptions_and_limitations_to_copyright.2C_such_as_fair_dealing_and_fair_use.3F">Mer information</a>.</p>
</div>
</div>
<div id="help_publicity_privacy_or_moral_rights_popup" class="help_panel">
<div class="bd">
<p>Du behöver få ytterligare tillstånd innan du använder materialet som du tänkt dig. </p>
<p><a href="https://wiki.creativecommons.org/Considerations_for_licensors_and_licensees">Mer information</a>.</p>
</div>
</div>
</div>
<script type='text/javascript' src='/wp-content/themes/cc/js/cc.js'></script>
<script type='text/javascript' src='/wp-content/plugins/cc-donate/js/cc-donate.js'></script>
<script type='text/javascript' src='/wp-content/themes/cc/js/breakpoint-body-class.js'></script>
<script type='text/javascript' src='/wp-content/themes/cc/js/sticky-nav.js'></script>
<script type='text/javascript' src='/wp-content/themes/cc/js/toggle-search.js'></script>
<script type='text/javascript' src='/wp-content/themes/cc/js/donation.js'></script>
<script type='text/javascript' src='/wp-content/themes/twentysixteen/js/skip-link-focus-fix.js'></script>
<script type='text/javascript'>
  /* <![CDATA[ */
  var screenReaderText = {"expand":"visa undermeny","collapse":"dölj undermeny"};
  /* ]]> */
  </script>
<script type='text/javascript' src='/wp-content/themes/twentysixteen/js/functions.js'></script>
<script type="text/javascript">
    //<![CDATA[
    var donateForms = $('.deed-donate-form');

    $(donateForms).each(function() {
      var otherFields = $('input[value="gf_other_choice"]');

      $(this).on('submit', function() {
        $(otherFields).each(function() {
          var parent = $(this).closest('li');
          var radioField = $(this);
          var txtField = $(parent).children('input[type="text"]');
          var txtValue = txtField.val();

          if (txtValue || radioField.is(':checked')) {
            radioField.val(txtValue);
          }
        });
      });
    });
    //]]>
  </script>
<script type="text/javascript">
    //<![CDATA[
    $(document).ready(function() {
        $('#deed-donate-slide').addClass('slider');
        $('#deed-donate-slide').show();
        // Set banner to reveal after X seconds
        setTimeout(function(){
            $('#deed-donate-slide').addClass('reveal');
        }, 5000);
        $(window).scroll(function() {
            if ($(window).scrollTop() <= 160) {
                $('#deed-donate-slide').finish();
                //$('#deed-donate-slide').removeClass('reveal');
            } else {
                $('#deed-donate-slide').addClass('reveal');
            }
        });

        $('.slide-close').click(function(event) {
            $('#deed-donate-slide').remove();
        });

        /* Close slider on pressing ESC */
        $(document).keyup(function(e) {
            if (e.keyCode === 27) {
                $('#deed-donate-slide').remove();
            }
        });

        $(".slide-trigger p, .slide-trigger button").click(function(){
            window.location.href = "https://us.netdonor.net/page/6650/donate/1?ea.tracking.id=deed-overlay";

        });
    });
    //]]>
  </script>
<script type="text/javascript">
    //<![CDATA[
    var _gaq = _gaq || [];
    _gaq.push(['_setAccount', 'UA-2010376-1']);
    _gaq.push(['_trackPageview']);
  
    (function() {
      var ga = document.createElement('script'); ga.type = 'text/javascript'; ga.async = true;
      ga.src = ('https:' == document.location.protocol ? 'https://ssl' : 'http://www') + '.google-analytics.com/ga.js';
      var s = document.getElementsByTagName('script')[0]; s.parentNode.insertBefore(ga, s);
    })();
    //]]>
  </script>

<script type="text/javascript">
    (function(w,d,s,l,i){w[l]=w[l]||[];w[l].push({'gtm.start':
    new Date().getTime(),event:'gtm.js'});var f=d.getElementsByTagName(s)[0],
    j=d.createElement(s),dl=l!='dataLayer'?'&l='+l:'';j.async=true;j.src=
    'https://www.googletagmanager.com/gtm.js?id='+i+dl;f.parentNode.insertBefore(j,f);
    })(window,document,'script','dataLayer','GTM-KP4CRCM');
  </script>


<noscript><iframe src="https://www.googletagmanager.com/ns.html?id=GTM-KP4CRCM"
  height="0" width="0" style="display:none;visibility:hidden"></iframe></noscript>

<script type="text/javascript">
    //<![CDATA[
    $(document).ready(function() {
      $('#deed .helpLink').each(function(index, helpLinkElem) {
        var helpId = $(helpLinkElem).attr('id');
        var popupId = helpId ? 'help_' + helpId : undefined;
        $(this).attr('tabindex',0);
        if (popupId) {
          var popupElem = $('#'+popupId);
          var popupTitleHtml = $('.hd', popupElem).html();
          var popupBodyHtml = $('.bd', popupElem).html();
          $(helpLinkElem).popover({
            placement: 'auto top',
            viewport: '#deed',
            trigger: 'focus',
            title: popupTitleHtml ? popupTitleHtml : undefined,
            content: popupBodyHtml ? popupBodyHtml : undefined,
            html: true
          });
        }
      });

      $('.helpLink').on('click', function(e) {
        e.preventDefault();
      });
    });
    //]]>
  </script>
<script type="text/javascript" src="/includes/language-selector.js"></script>
</body>
</html>